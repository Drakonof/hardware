`define MAC_WIDTH        48
`define IP_V4_WIDTH      32
`define UDP_WIDTH        16